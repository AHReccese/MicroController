`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:35:09 03/05/2019 
// Design Name: 
// Module Name:    FP_Pre2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 

//
//////////////////////////////////////////////////////////////////////////////////
module FP_Pre2(input[26:0] a,input [5:0]b ,output sticky_bit,output [26:0] result
    );
		
assign result[26:0] = a>>b[5:0];

assign sticky_bit =   							( b == 1 ) ? a[0] :
 							( b == 2 ) ? a[0]|a[1] :
 							( b == 3 ) ? a[0]|a[1]|a[2] :
 							( b == 4 ) ? a[0]|a[1]|a[2]|a[3] :
 							( b == 5 ) ? a[0]|a[1]|a[2]|a[3]|a[4]:
 							( b == 6 ) ? a[0]|a[1]|a[2]|a[3]|a[4]|a[5] :
 							( b == 7 ) ? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6] :
 							( b == 8 ) ? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7] :
 							( b == 9 ) ? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8] :
 							( b == 10) ? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9] :
 							( b == 11) ? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10] :
 							( b == 12 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11] :
 							( b == 13 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12] :
 							( b == 14 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13] :
 							( b == 15 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14] :
 							( b == 16 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15] :
 							( b == 17 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16] :
 							( b == 18 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17] :
 							( b == 19 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18] :
 							( b == 20 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19] :
 							( b == 21 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20] :
 							( b == 22 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21] :
 							( b == 23 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22] :
 							( b == 24 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23] :
 							( b == 25 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24] :
 							( b == 26 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25] :
 							( b == 27 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25]|a[26] :
 							( b == 28 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25]|a[26] :
 							( b == 29 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25]|a[26] :
 							( b == 30 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25]|a[26] :
 							( b == 31 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25]|a[26] :
 							( b == 32 )? a[0]|a[1]|a[2]|a[3]|a[4]|a[5]|a[6]|a[7]|a[8]|a[9]|a[10]|a[11]|a[12]|a[13]|a[14]|a[15]|a[16]|a[17]|a[18]|a[19]|a[20]|a[21]|a[22]|a[23]|a[24]|a[25]|a[26] : 0;
 								
endmodule
